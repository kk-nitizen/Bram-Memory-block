package datatypes;
import FixedPoint::*;
typedef FixedPoint#(16,16) DataType;
typedef UInt#(16) ImgWidth;
typedef FixedPoint#(2,14) CoeffType;
typedef UInt#(12) BramWidth;
typedef UInt#(6) BramLength;

endpackage
